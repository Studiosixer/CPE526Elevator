architecture behavioral of elevator is
begin

end architecture;